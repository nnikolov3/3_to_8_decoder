/*******************************************
Nikolay Nikolov
Project 1 Problem 2
Module of a 3 to 8 Decoder 
*******************************************/

//******************************************
module decoder (A,B,C,en,d0,d1,d2,d3,d4,d5,d6,d7);
//******************************************  
 output d0,d1,d2,d3,d4,d5,d6,d7;
 input A,B,C;
 input en;
  
  assign {d0, d1, d2, d3, d4, d5, d6, d7} = 
 ( {en,A,B,C} == 4'b1000) ? 8'b1000_0000 :
 ( {en,A,B,C} == 4'b1100) ? 8'b0100_0000 :
 ( {en,A,B,C} == 4'b1010) ? 8'b0010_0000 :
 ( {en,A,B,C} == 4'b1110) ? 8'b0001_0000 :
 ( {en,A,B,C} == 4'b1001) ? 8'b0000_1000 :
 ( {en,A,B,C} == 4'b1101) ? 8'b0000_0100 :
 ( {en,A,B,C} == 4'b1011) ? 8'b0000_0010 :
 ( {en,A,B,C} == 4'b1111) ? 8'b0000_0001 :
  8'b0000_0000;
  
endmodule